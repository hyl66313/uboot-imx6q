module
endmodule

